* DRIVER

.include ../BC547B.model
.include ../ponteh.model

VCC 10 0 DC 9
VIN1 20 0 PULSE(0 5 2NS 2NS 2NS 10MS 20MS)

R1 10 2 1000
Q1 2 20 0 BC547B
*C1 20 2 20p

* vcc ref v1+ v1- v2+ v2- vo+ vo-
xp1 10 0 20 2  5 6 ponteh

Rl 5 6 1000

* ANALYSIS
.TRAN 	.001S  .02S
*.AC 	DEC 	5 .1Hz 10000KHz
*

.control
 run
 plot   v(5) - v(6)
.endc



