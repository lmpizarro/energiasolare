POTENTIOSTAT.CIR
*
.include ../models/generics/diffStage.model


* POWER SUPPLIES
VCC	11	0	DC	+15
VDD	12	0	DC	-15

* SIGNAL SOURCE
*V60	1	0	SIN(0	1V	1KHZ)   AC
*V60 1 0  PULSE(500MV -500MV 0 0.000001 0.000001 0.005 .01)
V60 1 0  PULSE(-500MV 500MV 10NS 10NS 10NS 0.0005 .001)
*V60	1	0	DC       .001	

* Vcc Vdd v+ v- o+ o- 
xp1 11 12 1 0 5 6  diffStage 

C1 5 7 .1U
RL 7 0 100000



* ANALYSIS
.TRAN .001m 10mm
.AC 	DEC 	5 10Hz 10KHz
.PLOT	AC 	VM(7)
*

.control
run
 plot   v(7)  
.endc



