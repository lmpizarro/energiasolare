DOA1PNP.CIR
*
.include ../models/generics/doa1pnp.model
.include ../models/ci/ne5534.model


* POWER SUPPLIES
VCC	11	0	DC	+24
VDD	12	0	DC	-24

* SIGNAL SOURCE
V60	10	0	AC SIN(0	.060V	1KHZ)
*V60 1 0  PULSE(500MV -500MV 0 0.000001 0.000001 0.005 .01)
*V60 1 0  PULSE(-500MV 500MV 10NS 10NS 10NS 0.005 .01)
*V60	1	0	DC       0	


Rg 10 1 60000
* v+ v- Vcc Vdd  o 
xp1 1 8 11 12 7   doa1PNP 

RF1 7 8 60000
RF2 8 100 3000
C2 100 0 100u
*CF1 7 8 20p

C1 7 9 100u
Rl 9 0 600

* ANALYSIS
.TRAN .01m 10MS
.AC 	DEC 	10 1Hz 10000KHz
.PLOT	AC 	VM(7)
*

.control
run
 plot v(9) 
 *plot v(7)
 AC 	DEC 	10 1Hz 100000KHz
 plot vdb(9) 
.endc



