POTENTIOSTAT.CIR
*
.include ../models/generics/potentiostat.model


* POWER SUPPLIES
VCC	11	0	DC	+15
VDD	12	0	DC	-15

* SIGNAL SOURCE
*V60	1	0	SIN(0	1MVPEAK	100HZ)   AC
*V60 1 0  PULSE(500MV -500MV 0 0.000001 0.000001 0.0005 .001)
V60 1 0  PULSE(0MV 500MV 1uS 1uS 1uS 0.0005 1)
*V60	1	0	DC       .001	

* sig ref CE RE WE OUT
xp1 1 0 3 5 6 7 potentiostat

* randless
R4 3 5 2000K
R5 9 5 2000000
R6 9 6 100000 
C1 9 6 100u


* ANALYSIS
.TRAN .001m 1mm
.AC 	DEC 	5 .1Hz 100000KHz
.PLOT	AC 	VM(4)
*

.control
run
 plot   v(7) 
.endc



