j-918-clone.CIR 

.include ../models/generics/compounds.model
.include ../models/components/BC547B.model
.include ../models/components/BC557.model
.include ../models/generics/currSource.model
.include ../models/components/1n4148.model
.include ../models/components/TIP110.SP2
.include ../models/components/TIP117.SP3

*
* INPUT VOLTAGE
VCC	12	0	DC	15 
*sin(0v .01VPEAK 50HZ)
VDD	11	0	DC	-15
Vin1	1	0	AC  SIN(0  0.001VPEAK  1.0KHZ)
*Vin2	2	0	AC  SIN(0  -0.0VPEAK  1.0KHZ)

XO1 12 11 1 0 3 j918B
*XOU 12 11 1 3 OUTB

Rl 3 0 100000

.SUBCKT j918B 12 11 1 2 22 
D1 12 101 1N4148
D2 101 Bq3 1N4148
R7 Bq3 11 27000

r1 12 9 1300
q3 3 Bq3 9 BC557

re1 3 30 100
re2 3 31 100

q1 4 1 30 BC557
q2 5 2 31 BC557

rc1 4 11 8200

* CS q2
*r6 12 bq4 27000
*D3 bq4 8 1N4148
*D4 8 11 1N4148
*qc2 5 bq4 6 BC547B
*R5 6 11 2700

RC2 5 11 8200

Xout 12 11 5 22 OUTA

.ENDS j918B

.SUBCKT OUTa 12 11 5 22
RC 12 22 5000
XT1 22 5 23 Xtip110
RE 23 11 1
.ENDS OUTa

.SUBCKT OUTC 12 11 5 22
D5 12 13 1N4148
D6 13 14 1N4148
R8 14 11 27000
r9 12 15 150
xQ5 16 14 15 tip117

D7 16 17 1N4148
D8 17 18 1N4148

XT1 18 5 23 Xtip110
R2 23 11 150
C1 16 18 0.001u

D10 18 22 1N4148
D9 22 16 1N4148


.ENDS OUTC

.SUBCKT OUTB 12 11 5 22


D5 12 13 1N4148
D6 13 14 1N4148
R8 14 11 27000

r9 12 15 150
Q5 16 14 15 BC557

D7 16 17 1N4148
D8 17 18 1N4148
Q6 18 5 20 BC547B

R10 20 11 10000

Q7 18 20 21 BC547B
R11 21 11 150
C2 16 18 .001u
C1 18 19 36p
R12 19 5 470

D10 18 22 1N4148
D9 22 16 1N4148

q8 11 16 23 BC547B
R14 23 22 4.7

q9 11 18 24 BC557
R13 24 22 4.7


.ENDS OUTB

.SUBCKT j918 12 11 1 2 16

XCS1 12 11 7 CURRSRCPNP RI = 1300 RB = 17000

*XCS2 12 11 16 CURRSRCNPN RI = 270 RB = 17000


Re1 7 13 100
Re2 7 14 100

XSZ1 9 1 13 SZKPNP
XSZ2 16 2 14 SZKPNP

RC2 16 11 8200
RC1 9 11 8200

.ENDS j918

*
* ANALYSIS
.TRAN 	0.001MS  	10.0MS
.ac dec 10 1 10MHZ
*.disto 	dec 10 20 20000
*.noise v(8) vin dec 10 1 2000000
*
.control
run
plot v(3)
ac dec 10 1 100000000
plot vdb(3)
.endc

* VIEW RESULTS
.PRINT	TRAN V(8) 
.PROBE
.END
