DIFFSTAGEPNP.CIR
*
.include ../models/generics/diffStageSZP.model
.include ../models/generics/opamp1.model
.include ../models/ci/ne5534.model


* POWER SUPPLIES
VCC	11	0	DC	+15
VDD	12	0	DC	-15

* SIGNAL SOURCE
V60	1	0	SIN(0	.3V	1KHZ)   AC
*V60 1 0  PULSE(500MV -500MV 0 0.000001 0.000001 0.005 .01)
*V60 1 0  PULSE(-500MV 500MV 10NS 10NS 10NS 0.0005 .001)
*V60	1	0	DC       .001	

* Vcc Vdd v+ v- o+ o- 
xp1 11 12 1 0 5 6  diffStageSZP 

xopamp1 6 7 7 opamp1 
xopamp2 5 8 8 opamp1 

R3 7 10 10000
R2 15 10 11000
R4 8 9 10000
R5 9 0 11000

Xopamp3 9 10 15 opamp1



* ANALYSIS
.TRAN .01m 2mm
.AC 	DEC 	5 10Hz 10KHz
.PLOT	AC 	VM(7)
*

.control
run
 plot     v(15)
 *plot v(7) 
 *plot v(5) - v(6) xlimit 0.0004995 0.0005005
.endc



