* DRIVER

.include ../models/BC547B.model
.include ../models/BC557.model
.include ../models/sihf630.lib
.include ../models/sihf540.lib
.include ../models/irf530.lib
.include ../models/irf510.lib
.incude ../models/1N4148B.model
.incude ../models/TIP110.SP3
.include ../models/TIP31.SP3
.include ../models/bav21.model

VCC 10 0 DC 9
VIN1 20 0 PULSE(0 9V 1NS 1NS 1NS .005MS .01MS)

*D1 20 1  1N4148B
RP 1 0 1000
L1 10 2 200u
Q1 0 20 1 BC557
XQ1 2 1 0 irf510
Q2 10 20 1 BC547B

D2 2 3 bav21

Cl 3 0 100u
Rl 3 0 10000


* ANALYSIS
.TRAN 	.00001S  .00005S
*.AC 	DEC 	5 .1Hz 10000KHz
*

.control
 run
 plot   v(2)
.endc



