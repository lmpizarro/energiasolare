CURRENTsOURCE.CIR

.include ../models/components/BD140B.LIB
.include ../models/components/BD139.SP3
.include ../models/components/1n4148.model


* INPUT VOLTAGE
VCC	11	0	DC	25 
VDD	12	0	DC	-25
Vin1	1	0	AC  SIN(0  0.100100VPEAK  1.0KHZ)


RIN 1 100 150


RS 11 10 1.2K
q1 9 10 11 bc560C
RP 9 12 30K
q2 3 9 10 bc560C

q3 800 nf2 3 BC560C
q4 600 100 3 BC560C

qs3 3 800 8 bc550C
qs4 3 600 6 bc550C
rski1 800 8 10K
rski2 600 6 10K


q5 6 8 7 bc550C
q6 8 7 12 bc550C
q7 7 7 12 bc550C


* ---------------  Output ---------------
*RC1 11 16 10K

RC1 11 165 130
RC1P 164 12 10K
Q202 16 164 165 BC560C
Q201 164 165 11 BC560C


q10 16 16 15 bc550C
q11 15 15 14 bc550C 

RSK 14 13 1.0K
q8 13 6 120 bc550C
q9 120 13 14 bc560C
resk 120 12 200


q12 31 16 17 bc550C 
Q13 32 14 19 bc560C
re5 17 18 4.7
re6 18 19 4.7
res5 31 11 500
res6 32 12 500

q14 17 31 11 BC327
q15 19 32 12 BC337

rf1 18 nf2 10K
**cf1 18 nf2 90p
rf2 nf2 20 100
CP 20 0 500u

ccp 60 6 40p
rcp 60 14 300

RL 18 0 600


.SUBCKT ICM_N 1 2 3
* VCC VDD out
R1 1 4 30K
RS 5 2 1.2K
Q1 4 5 2 bc547a
Q2 3 4 5 bc547a 
.ENDS

.SUBCKT ICM_P 1 2 3
* VDD VCC out

R1 1 4 10K
RS 5 2 .1K
Q1 4 5 2 bc557a
Q2 3 4 5 bc557a 

.ENDS

.SUBCKT IDIFF 1 2 3
* IN VDD  out

Q1 1 4 2 bc547a 
Q2 4 4 2 bc547a
Q3 3 1 4 bc547a 
.ENDS 

.SUBCKT DIFF 1 2 3 4 5
* V- V+ CM 4 out

RE1 3 5 20
RE2 3 6 20

XQ1 4 1 5 BD140
XQ2 5 2 6 BD140

.ENDS

.SUBCKT OFFCMP 1 3 4 0
* VCC in+ in- ref
R1 1 2 5K
R2 2 0 5K

r3 5 2 1M
r4 6 2 1M
r5 3 5 1M
r6 4 6 1N
c1 5 0 1u
c2 6 0 1u
.ENDS

.model bc547a NPN BF=400 NE=1.3 ISE=10.3F IKF=50M IS=10F VAF=80 ikr=12m
       + BR=9.5 NC=2 VAR=10 RB=280 RE=1 RC=40 VJE=.48 tr=.3u tf=.53n
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47p kf=2f
.model bc547b NPN BF=500 NE=1.3 ISE=9.72F IKF=80M IS=20F VAF=50 ikr=12m
       + BR=10 NC=2 VAR=10 RB=280 RE=1 RC=40 VJE=.48 tr=.3u tf=.53n
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47p kf=2f
.model bc547c NPN BF=730 NE=1.4 ISE=29.5F IKF=80M IS=60F VAF=25 ikr=12m
       + BR=10 NC=2 VAR=10 RB=280 RE=1 RC=40 VJE=.48 tr=.3u tf=.53n
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47.6p kf=2f
.model BC557a PNP BF=190 NE=1.5 ISE=12F IKF=90M IS=10F VAF=50 ikr=12m
       + nc=2 br=4 var=10 rb=280 re=1 rc=40 vje=.48 tf=.5n tr=.3u
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47.6p kf=2f
.model BC557b PNP BF=335 NE=1.5 ISE=7.35F IKF=82M IS=10F VAF=40 ikr=12m
       + nc=2 br=4 var=10 rb=280 re=1 rc=40 vje=.48 tf=.5n tr=.3u
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47.6p kf=2f
.model BC557c PNP BF=490 NE=1.5 ISE=12.4F IKF=78M IS=60F VAF=36 ikr=12m
       + nc=2 br=4 var=10 rb=280 re=1 rc=40 vje=.48 tf=.5n tr=.3u
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47.6p kf=2f
.model BD140 pnp IS=1e-09 BF=650.842 NF=0.85 VAF=10 IKF=0.0950125 ISE=1e-08 NE=1.54571 
       +BR=56.177 NR=1.5 VAR=2.11267 IKR=0.950125 ISC=1e-08 NC=3.58527 RB=41.7566 
       +IRB=0.1 RBM=0.108893 RE=0.000347052 RC=1.32566 XTB=19.5239 XTI=1 EG=1.05 
       +CJE=1e-11 VJE=0.75 MJE=0.33 TF=1e-09 XTF=1 VTF=10 ITF=0.01
       +CJC=1e-11 VJC=0.75 MJC=0.33 XCJC=0.9 FC=0.5 CJS=0 VJS=0.75 
       +MJS=0.5 TR=1e-07 PTF=0 KF=0 AF=1
.MODEL Qbd136 pnp IS=1e-09 BF=681.414 NF=0.85 VAF=10 IKF=0.196957 ISE=1e-08 NE=1.57381 
       +BR=56.5761 NR=1.5 VAR=0.975138 IKR=0.952908 ISC=1e-08 NC=3.58666 RB=40.4245 
       +IRB=0.1 RBM=0.106663 RE=0.00034585 RC=1.31191 XTB=22.4074 XTI=1 EG=1.05 
       +CJE=1e-11 VJE=0.75 MJE=0.33 TF=1e-09 XTF=1 VTF=10 ITF=0.01
       +CJC=1e-11 VJC=0.75 MJC=0.33 XCJC=0.9 FC=0.5 CJS=0 VJS=0.75 MJS=0.5
       +TR=1e-07 PTF=0 KF=0 AF=1
.MODEL BC550C npn IS=45e-15 BF=689 VAF=162 IKF=0.09 ISE=4600e-15 NE=1622 NF=0.9965
       +RB=167 RC=1RE=0.04 CJE=18.7e-12 MJE=0.35 VJE=0.75
       +CIRJC=6.2e-12 MJC=0.25 VJC=0.4 FC=0.5
       +TF=595e-12 XTF=10 VTF=10 ITF=15NE TR=10e-9 BR=12.2 IKR=0.34
       +EG=1.2 XTB=1.65 XTI=3 NC=0.996 NR=1.08 VAR=120 IRB=7e-5 RBM=1.1
       +XCJC=0.6 ISC=5e-15
.MODEL BC560C pnp IS=60e-15 BF=300 VAF=160
       +IKF=0.10 ISE=70e-15 NE=1.42 NF=1 RB=170	RC=1.0	RE=0.05
       +CJE=19e-12 MJE=0.3 VJE=0.75 CJC=3.9e-12	MJC=0.3	VJC=0.75 FC=0.5
       +TF=600e-12 XTF=7 VTF=4	ITF=0.45 TR=10e-9 BR=3	IKR=0
       +EG=1.1 XTB=1.5 XTI=3 NC=2 ISC=0	
.MODEL BD139C npn
+IS=150e-15	BF=260 		VAF=99
+IKF=1.2	ISE=70e-15	NE=1.2		NF=1.0
+RB=5		RC=0.01		RE=0.08
+CJE=293e-12 	MJE=0.33	VJE=0.67
+CJC=49e-12	MJC=0.39	VJC=0.52	FC=0.5
+TF=585e-12 	XTF=10000	VTF=35		ITF=20
+TR=10e-9	BR=78		IKR=0.14
+EG=1.21 	XTB=1.14	XTI=3		NC=1.45
+ISC=19e-12	NR=1.0		VAR=7.5		IRB=0.03
+RBM=0.001	XCJC=0.53
.MODEL BD140C pnp
+IS=120e-15	BF=113 		VAF=140
+IKF=1.5	ISE=1000e-15	NE=1.5		NF=1
+RB=5		RC=0.01		RE=0.1
+CJE=220e-12 	MJE=0.35	VJE=0.7
+CJC=68e-12	MJC=0.35	VJC=0.6		XCJC=0.5	FC=0.5
+TF=320e-12 	XTF=10000 	VTF=35		ITF=20
+TR=100e-9	BR=25		IKR=0.1		
+EG=1.2 	XTB=1.5		XTI=3		NC=1.4
+ISC=7e-12	NR=1.0		VAR=8		IRB=0.01	RBM=0.01	
.model BC327 PNP IS=1.08E-13 NF=0.99 ISE=2.713E-14 NE=1.4 BF=385.7 IKF=0.3603 
+VAF=31.29 NR=0.9849 ISC=5.062E-13 NC=1.295 BR=20.57 IKR=0.054 VAR=11.62 
+RB=1 IRB=1.00E-06 RBM=0.5 RE=0.1415 RC=0.2623 XTB=0 EG=1.11 XTI=3 
+CJE=5.114E-11 VJE=0.8911 MJE=0.4417 TF=7.359E-10 XTF=1.859 VTF=3.813 ITF=0.4393 
+PTF=0 CJC=2.656E-11 VJC=0.62 MJC=0.4836 XCJC=0.459 TR=5.00E-08 CJS=0 
+VJS=0.75 MJS=0.333 FC=0.99 Vceo=45 
.model BC337 NPN IS=4.13E-14 NF=0.9822 ISE=3.534E-15 NE=1.35 BF=292.4 IKF=0.9 
+VAF=145.7 NR=0.982 ISC=1.957E-13 NC=1.3 BR=23.68 IKR=0.1 VAR=20 RB=60 IRB=2.00E-04 
+RBM=8 RE=0.1129 RC=0.25 XTB=0 EG=1.11 XTI=3 CJE=3.799E-11 VJE=0.6752 
+MJE=0.3488 TF=5.4E-10 XTF=4 VTF=4.448 ITF=0.665 PTF=90 CJC=1.355E-11 
+VJC=0.3523 MJC=0.3831 XCJC=0.455 TR=3.00E-08 CJS=0 VJS=0.75 MJS=0.333 
+FC=0.643 Vceo=45 





.TRAN 	0.001MS  	10.0MS
.ac dec 10 1 10MHZ
.control
run
plot i(Vin1)  
plot v(18)
ac dec 10 1 100000000
plot vdb(18)
.endc


