POTENTIOSTAT.CIR
*
.include ../models/generics/potentiostat.model


* POWER SUPPLIES
VCC	11	0	DC	+15
VDD	12	0	DC	-15

* SIGNAL SOURCE
*V60	1	0	SIN(0	1MVPEAK	100HZ)   AC
*V60 1 0  PULSE(500MV -500MV 0 0.000001 0.000001 0.005 .01)
V60 1 0  PULSE(0MV 500MV 10NS 10NS 10NS 0.005 1)
*V60	1	0	DC       .001	

* sig ref CE RE WE OUT
xp1 1 0 3 5 6 7 potentiostat

* randless
R4 3 5 20K
R5 5 9 10000
R6 9 6 100000 
C1 9 6 1u


* ANALYSIS
.TRAN .001m 50mm
.AC 	DEC 	5 10Hz 10KHz
.PLOT	AC 	VM(7)
*

.control
run
 plot   v(7) 
.endc



