* TESTIRF630
* info: https://threeneurons.wordpress.com/nixie-power-supply/hv-supply-kit/

.include ../models/components/BC547B.model
.include ../models/components/BC557.model
.include ../models/components/sihf630.lib
.include ../models/components/sihf540.lib
.include ../models/components/irf530.lib
.include ../models/components/irf510.lib
.incude ../models/components/1N4148B.model
.incude ../models/components/TIP110.SP3
.include ../models/components/TIP31.SP3
.include ../models/components/bav21.model

VCC 10 0 DC 9
VIN1 20 0 PULSE(0 9V 1NS 1NS 1NS .005MS .01MS)

*D1 20 1  1N4148B
RP 1 0 1000
L1 10 2 200u
Q1 0 20 1 BC557
XQ1 2 1 0 irf510
Q2 10 20 1 BC547B

D2 2 3 bav21

Cl 3 0 100u
Rl 3 0 10000


* ANALYSIS
.TRAN 	.00001S  .00005S
*.AC 	DEC 	5 .1Hz 10000KHz
*

.control
 run
 plot   v(2)
.endc



