CURRENTsOURCE.CIR

.include ../models/components/BD140B.LIB
.include ../models/components/BD139.SP3
.include ../models/components/1n4148.model


* INPUT VOLTAGE
VCC	11	0	DC	25 
VDD	12	0	DC	-25
Vin1	1	0	AC  SIN(0  0.100100VPEAK  1.0KHZ)


RIN 1 100 150


RS 11 10 1.2K
q1 9 10 11 bc557a
RP 9 12 30K
q2 3 9 10 bc557a


q3 8 nf2 3 QBD140
q4 6 100 3 QBD140

q5 6 8 7 bc547a
q6 8 7 12 bc547a
q7 7 7 12 bc547a


*RC1 11 16 10K

RC1 11 165 135
RC1P 164 12 10K
Q202 16 164 165 BC557a
Q201 164 165 11 BC557a


q10 16 16 15 bc547a
q11 15 15 14 bc547a 

RSK 14 13 1.0K
q8 13 6 120 bc547a
q9 120 13 14 bc557a
resk 120 12 200

*q8 14 6 12 bc547a

q12 11 16 17 bc547a 
Q13 12 14 19 bc557a
re5 17 18 4.7
re6 18 19 4.7

rf1 18 nf2 50K
**cf1 18 nf2 90p
rf2 nf2 20 100
CP 20 0 500u

ccp 60 6 40p
rcp 60 14 300


.SUBCKT ICM_N 1 2 3
* VCC VDD out
R1 1 4 30K
RS 5 2 1.2K
Q1 4 5 2 bc547a
Q2 3 4 5 bc547a 
.ENDS

.SUBCKT ICM_P 1 2 3
* VDD VCC out

R1 1 4 10K
RS 5 2 .1K
Q1 4 5 2 bc557a
Q2 3 4 5 bc557a 

.ENDS

.SUBCKT IDIFF 1 2 3
* IN VDD  out

Q1 1 4 2 bc547a 
Q2 4 4 2 bc547a
Q3 3 1 4 bc547a 
.ENDS 

.SUBCKT DIFF 1 2 3 4 5
* V- V+ CM 4 out

RE1 3 5 20
RE2 3 6 20

XQ1 4 1 5 BD140
XQ2 5 2 6 BD140

.ENDS

.SUBCKT OFFCMP 1 3 4 0
* VCC in+ in- ref
R1 1 2 5K
R2 2 0 5K

r3 5 2 1M
r4 6 2 1M
r5 3 5 1M
r6 4 6 1N
c1 5 0 1u
c2 6 0 1u
.ENDS

.model bc547a NPN BF=400 NE=1.3 ISE=10.3F IKF=50M IS=10F VAF=80 ikr=12m
       + BR=9.5 NC=2 VAR=10 RB=280 RE=1 RC=40 VJE=.48 tr=.3u tf=.5n
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47p kf=2f
.model bc547b NPN BF=500 NE=1.3 ISE=9.72F IKF=80M IS=20F VAF=50 ikr=12m
       + BR=10 NC=2 VAR=10 RB=280 RE=1 RC=40 VJE=.48 tr=.3u tf=.5n
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47p kf=2f
.model bc547c NPN BF=730 NE=1.4 ISE=29.5F IKF=80M IS=60F VAF=25 ikr=12m
       + BR=10 NC=2 VAR=10 RB=280 RE=1 RC=40 VJE=.48 tr=.3u tf=.5n
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47.6p kf=2f
.model BC557a PNP BF=190 NE=1.5 ISE=12F IKF=90M IS=10F VAF=50 ikr=12m
       + nc=2 br=4 var=10 rb=280 re=1 rc=40 vje=.48 tf=.5n tr=.3u
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47.6p kf=2f
.model BC557b PNP BF=335 NE=1.5 ISE=7.35F IKF=82M IS=10F VAF=40 ikr=12m
       + nc=2 br=4 var=10 rb=280 re=1 rc=40 vje=.48 tf=.5n tr=.3u
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47.6p kf=2f
.model BC557c PNP BF=490 NE=1.5 ISE=12.4F IKF=78M IS=60F VAF=36 ikr=12m
       + nc=2 br=4 var=10 rb=280 re=1 rc=40 vje=.48 tf=.5n tr=.3u
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc:.33 isc=47.6p kf=2f



.TRAN 	0.001MS  	10.0MS
.ac dec 10 1 10MHZ
.control
run
plot i(Vin1)  
plot v(18)
ac dec 10 1 100000000
plot vdb(18)
.endc


