* HWRSPLIT

.include ../models/generics/doubler.model

VIN1 80 0 ac 1.0 sin(0.0 33.84 50.0 0 0)

* vi 0 v+ v- 
xp1 80 0 5   doubler

Rl1 5 0 5000


* ANALYSIS
.TRAN 	.001S  2S
*.AC 	DEC 	5 .1Hz 10000KHz
*

.control
 run
 plot    v(5)
.endc



