BASIC_AMPLIFIER.CIR - DISCRETE AMPLIFIER
*
.include ../components/1n4148w.txt
.include ../components/BC547B.SP3
.include ../components/BC557B.SP3
.include ../components/bd139.lib
.include ../components/bd140.lib

*
* POWER SUPPLIES
VCC	100	0	DC	+25V
VEE	101	0	DC	-25V


VS	1	0	AC 1	SIN(0 0.01V 1KHZ)
*CIN	1	2	1UF
*RIN1	2	0	100K


xop 100 101 1 3 20 opamp4

* FEEDBACK
RF2	20	3	33K
RF1	3	30	.15K
CF2     30  0 1000u
CCF1	20	3	5pF

* LOAD
RL	20	0	600

.subckt opamp4 100 101 2 3  20
* DIFF AMP

*xRECS	100	101 8 CURRSRCPNP RI = 1.3K	

xQ1	4 2 	8	SZKPNP
xQ2	40 3	8	SZKPNP

QC1 40 40 101 BC547B
QC2 4 40 101 BC547B

*RC1	4	101	1800
*XRCS1 100 101 4 CURRSRCNPN RI = 2600
*CC1	101	4	10PF
*
* GAIN STAGE AND COMPENSATION
XQ3	14 4	1010	SZKNPN
REq3 1010 101 150
CC2	14	4	270PF
*
* OUTPUT STAGE BIAS
*xRC3	100	101 11 CURRSRCPNP RI = 175	
xRCx2	100	101 8 11 CURRSRCx2PNP RI1 = 1.3K RI2 = 175	

xD1	11	13	D1N4148
xD2	13	14	D1N4148
*
* OUTPUT STAGE
Q4	100 11	200	QBD139
Q5	101 14	201	QBD140
RE1 200 20 10
RE2 201 20 10
*Qp1 11 200 20 BC547B
*Qp2 14 201 20 BC557B
DCl1 20 13 D1N4148
DCl2 13 20 D1N4148
*
*
.ENDS OPAMP4

.SUBCKT SZKNPN 1 2 3
q1 4 2 3 BC547B
q2 3 4 1 BC557B
R1 4 1 3K
C1 4 2 15p
.ENDS SZKPNP

.SUBCKT SZKPNP 1 2 3
q1 4 2 3 BC557B
q2 3 4 1 BC547B
R1 4 1 4K
.ENDS SZKPNP

.SUBCKT CURRSRCPNP 1 2 3  RI = 175 
Q1 3 4 5 BC557B
D1 1 6 D1N4148
D2 6 4 D1N4148
R1 4 2 24K
R2 5 1 {RI}
.ENDS CURRSRCPNP

.SUBCKT CURRSRCNPN 1 2 3  RI = 2700 
Q1 3 4 5 BC547B
D1 4 6 D1N4148
D2 6 2 D1N4148
R1 1 4 24K
R2 5 2 {RI}
.ENDS CURRSRCNPN

.SUBCKT CURRSRCx2PNP 1 2 3 7  RI1 = 175  RI2 = 150
Q1 3 4 5 BC557B
D1 1 6 D1N4148
D2 6 4 D1N4148
R1 4 2 24K
R2 5 1 {RI1}

Q2 7 4 8 BC557B

R3 8 1 {RI2}
.ENDS CURRSx2RCPNP


*
* SMALL SIGNAL DEVICES
.model	QNPN	NPN(BF=100)
.model	QPNP	PNP(BF=100)
.model	QNPN3	NPN(BF=100)
.model	D1N4148B	D(Is=0.1p Rs=16 CJO=2p Tt=12n Bv=100 Ibv=0.1p)

* OUTPUT POWER DEVICES
.model	QNPN4	NPN(BF=100)
.model	QPNP5	PNP(BF=100)

*
.TRAN	50US 20MS
.AC DEC 5 1 1MEG
.PROBE

.control
run
plot v(20) 
ac dec 10 1 100000000
plot vdb(20)
.endc
.END
