* test phvcell
.include ../models/generics/phvcell.model

X1 1 0 PHVCELL PARAMS: Iirr=4 


R1 1 0  100

* ANALYSIS
.TRAN 	.0001S  2S
*.AC 	DEC 	5 .1Hz 10000KHz
*

.control
 run
 plot  v(1)
.endc




